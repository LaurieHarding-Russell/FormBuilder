{
    "font" : "Bangers-Regular",
    "fontSize" : 100,
    "background": [1.0, 0, 0, 1.0],
    "height": "10%"
}