{
    "background" : [0.1, 0, 0.0, 1.0],
    "class1" : {
        "background" : [0.2, 0.0, 0.0, 1.0],
        "class2" : {
            "background" : [0.3, 0.0, 0.0, 1.0]
        }
    }
}