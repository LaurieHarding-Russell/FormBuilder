{
    background: [0.1, 0.5, 0.5, 0.5],
    class1 {
        background: [0.2, 0.5, 0.5, 0.5]
        class2 {
           background: [0.3, 0.5, 0.5, 0.5]
        }
    }
}