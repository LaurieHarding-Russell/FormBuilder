{
    "font" : "Bangers-Regular",
    "fontSize" : 100,
    "background": [1.0, 0, 0, 0.5],
    "width": "50%"
}