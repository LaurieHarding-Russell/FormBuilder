{
    "class1": {
        "height": "50%"
    }
}